
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY MO10 IS
END MO10;
 
ARCHITECTURE behavior OF MO10 IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT moshi
    PORT(
         CP : IN  std_logic;
         Rd : IN  std_logic;
         Q : OUT  std_logic_vector(3 downto 0);
         NQ : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal CP : std_logic := '0';
   signal Rd : std_logic := '0';

 	--Outputs
   signal Q : std_logic_vector(3 downto 0);
   signal NQ : std_logic_vector(3 downto 0);
   -- No clocks detected in port list. Replace CP below with 
   -- appropriate port name 
 
   constant CP_period : time := 60 ns;
 

BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: moshi PORT MAP (
          CP => CP,
          Rd => Rd,
          Q => Q,
          NQ => NQ
        );

   -- Clock process definitions
   CP_process :process
   begin
		CP <= '0';
		wait for CP_period/2;
		CP <= '1';
		wait for CP_period/2;
   end process;
 	

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
		 Rd<='0';
      wait for 100 ns;	
Rd<='1';
wait for CP_period*10;
		wait for CP_period*10;
		wait for CP_period*10;
		wait for CP_period*10;
		wait for CP_period*10;
      wait for CP_period*10;
wait for CP_period*10;
		wait for CP_period*10;
		wait for CP_period*10;
		wait for CP_period*10;
		wait for CP_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
